../vhdl_ecd_submodule/vhdl/spi_slave.vhd