../chisel/verilog/spi_slave.v