../vhdl_ecd_submodule/vhdl/synchronizer_n.vhd